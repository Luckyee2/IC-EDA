module acsoc04_1v8 ( EN, VDDA, VSSA, CS3_8u, CS2_4u, CS1_2u, CS0_1u );

  input CS2_4u;
  input CS0_1u;
  input EN;
  input VSSA;
  input VDDA;
  input CS1_2u;
  input CS3_8u;

  wire real CS0_1u;
  wire real CS0_2u;
  wire real CS0_4u;
  wire real CS0_8u;

  // Outputs declared as inputs so they can be tied together.
endmodule
